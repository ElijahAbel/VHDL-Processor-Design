library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity instructMem is
port (
  instructAddr : in std_logic_vector(31 downto 0); --input instruction from PC
  rd           : out std_logic_vector(31 downto 0) --output instruction to decoder and register file
);
end instructMem;

architecture rtl of instructMem is

-- --OPCODES
-- signal ARITH    : std_logic_vector(5 downto 0) := "000000"; --OPCODE00
-- signal ADDIMM   : std_logic_vector(5 downto 0) := "000001"; --OPCODE01
-- signal SUBIMM   : std_logic_vector(5 downto 0) := "000010"; --OPCODE02
-- signal ANDIMM   : std_logic_vector(5 downto 0) := "000011"; --OPCODE03
-- signal ORIMM    : std_logic_vector(5 downto 0) := "000100"; --OPCODE04
-- signal SHFLFT   : std_logic_vector(5 downto 0) := "000101"; --OPCODE05
-- signal LOAD     : std_logic_vector(5 downto 0) := "000111"; --OPCODE07
-- signal STORE    : std_logic_vector(5 downto 0) := "001000"; --OPCODE08
-- signal BLT      : std_logic_vector(5 downto 0) := "001001"; --OPCODE09
-- signal BEQ      : std_logic_vector(5 downto 0) := "001010"; --OPCODE0A
-- signal BNE      : std_logic_vector(5 downto 0) := "001011"; --OPCODE0B
-- signal JUMP     : std_logic_vector(5 downto 0) := "001100"; --OPCODE0C
-- signal HALT     : std_logic_vector(5 downto 0) := "111111"; --OPCODE3F

-- --FUNCTIONS
-- signal ADDREG   : std_logic_vector(5 downto 0) := "000001"; --FUNC1
-- signal SUBREG   : std_logic_vector(5 downto 0) := "000011"; --FUNC3
-- signal ANDREG   : std_logic_vector(5 downto 0) := "000101"; --FUNC5
-- signal ORREG    : std_logic_vector(5 downto 0) := "000111"; --FUNC7
-- signal NORREG   : std_logic_vector(5 downto 0) := "001001"; --FUNC9

begin

instruct : process (instructAddr)
begin
case instructAddr(31 downto 0) is
                            -- OPCODE&   RS    &  RT     &  RD     &  SHAMT  & FUNCT (R-TYPE)
				            -- OPCODE&   RS    &  RT     & Address/Immediate         (I-TYPE)
				            -- OPCODE&   Address (26-bits)                           (J-TYPE)
  when x"00000000" => rd <= "000111" & "00000" & "00010" & "00000" & "00000" & "011010";  --LB R2, R0, 26 //R2=A
  when x"00000004" => rd <= "000111" & "00000" & "00011" & "00000" & "00000" & "011011";  --LB R3, R0, 27 //R3=B
  when x"00000008" => rd <= "000001" & "00000" & "01001" & "00000" & "00000" & "001101";  --ADDI R9, R0, 13 //R9 to be used as the loop bound
  when x"0000000C" => rd <= "000111" & "00001" & "00100" & "00000" & "00000" & "000000";  --LB R4, R1, 0 //R4 holds S[i]
  when x"00000010" => rd <= "000111" & "00001" & "00101" & "00000" & "00000" & "000001";  --LB R5, R1, 1 //R5 holds S[i+1]
  when x"00000014" => rd <= "000000" & "00010" & "00100" & "00010" & "00000" & "000001";  --ADD R2, R2, R4
  when x"00000018" => rd <= "000000" & "00011" & "00101" & "00011" & "00000" & "000001";  --ADD R3, R3, R5
  when x"0000001C" => rd <= "000001" & "00001" & "00001" & "00000" & "00000" & "000001";  --ADDI R1, R1, 1 // R1 = 1 because 1 is the beginning value of i for our loop
  when x"00000020" => rd <= "000000" & "00010" & "00011" & "11100" & "00000" & "001001";  --NOR R28, R2 , R3  //R28 = A NOR B   --- Loop should come back to this line
  when x"00000024" => rd <= "000000" & "00010" & "11100" & "11101" & "00000" & "001001";  --NOR R29, R2 , R28 //R29 = A NOR R28
  when x"00000028" => rd <= "000000" & "00011" & "11100" & "11110" & "00000" & "001001";  --NOR R30, R3 , R28 //R30 = B NOR R28
  when x"0000002C" => rd <= "000000" & "11101" & "11110" & "11111" & "00000" & "001001";  --NOR R31, R29, R30 //R31 = R29 NOR R30
  when x"00000030" => rd <= "000000" & "11111" & "11111" & "00110" & "00000" & "001001";  --NOR R6 , R31, R31 //R6  = R31 NOR R31 (A XOR B)
  when x"00000034" => rd <= "000001" & "00110" & "01110" & "00000" & "00000" & "000000";  --ADDI R14,R6,0 //Store XOR value in R14
  when x"00000038" => rd <= "000011" & "00011" & "01010" & "00000" & "00000" & "011111";  --ANDI R10,R3,31 //Extracting 5 LSBs of B to find out the value to left rotate by, R11 contains the valu
  when x"0000003C" => rd <= "001010" & "01010" & "00000" & "00000" & "00000" & "000101";  --BEQ R10, R0, 5 //Skips SHL because R10 is 0
  when x"00000040" => rd <= "000001" & "00000" & "01011" & "00000" & "00000" & "000000";  --ADDI R11,R0,0 //Store 0 for our counter
  when x"00000044" => rd <= "000101" & "00110" & "00110" & "00000" & "00000" & "000001";  --SHL  R6 ,R6,1
  when x"00000048" => rd <= "000001" & "01011" & "01011" & "00000" & "00000" & "000001";  --ADDI R11, R11, 1 //increment R11
  when x"0000004C" => rd <= "001010" & "01010" & "01011" & "00000" & "00000" & "000001";  --BEQ, R10, R11, 1
  when x"00000050" => rd <= "001100" & "00000" & "00000" & "00000" & "00000" & "010001";  --JUMP 17
  when x"00000054" => rd <= "000001" & "00000" & "01100" & "00000" & "00000" & "100000";  --ADDI R12, R0, 32 //R12 = 32
  when x"00000058" => rd <= "000000" & "01100" & "01010" & "01100" & "00000" & "000011";  --SUB  R12, R12, R10 //R12 = 32 - LSB of B
  when x"0000005C" => rd <= "000001" & "00000" & "01101" & "00000" & "00000" & "000001";  --ADDI R13, R0, 1 //R13 = 1 if we are about to right shift A xor B
  when x"00000060" => rd <= "001100" & "00000" & "00000" & "00000" & "00000" & "111001";  --***CHANGED BY E**** JUMP 57 //after the halt
  when x"00000064" => rd <= "000000" & "00110" & "01110" & "00010" & "00000" & "000001";  --ADD R2, R6, R14 //Adding the left shifted and right shifted components together.
  when x"00000068" => rd <= "000101" & "00001" & "00111" & "00000" & "00000" & "000001";  --SHL R7, R1, 1 //R7 = 2xi
  when x"0000006C" => rd <= "000111" & "00111" & "01000" & "00000" & "00000" & "000000";  --LB R8, R7, 0 //R8 = S[2xi] 
  when x"00000070" => rd <= "000000" & "00010" & "01000" & "00010" & "00000" & "000001";  --ADD R2, R2, R8 //A = ((A xor B) << B) + S[2xi]
  when x"00000074" => rd <= "000000" & "00011" & "00010" & "11100" & "00000" & "001001";  --NOR R28, R3, R2 //R28 = B NOR A   --- Loop should come back to this line
  when x"00000078" => rd <= "000000" & "00011" & "11100" & "11101" & "00000" & "001001";  --NOR R29, R3, R28 //R29 = B NOR R28
  when x"0000007C" => rd <= "000000" & "00010" & "11100" & "11110" & "00000" & "001001";  --NOR R30, R2, R28 //R30 = A NOR R28
  when x"00000080" => rd <= "000000" & "11101" & "11110" & "11111" & "00000" & "001001";  --NOR R31, R29, R30 //R31 = R29 NOR R30
  when x"00000084" => rd <= "000000" & "11111" & "11111" & "00110" & "00000" & "001001";  --NOR R6, R31, R31 //R6 = R31 NOR R31 (B XOR A)
  when x"00000088" => rd <= "000001" & "00110" & "01110" & "00000" & "00000" & "000000";  --ADDI R14,R6,0 //Store XOR value in R14
  when x"0000008C" => rd <= "000011" & "00010" & "01010" & "00000" & "00000" & "011111";  --ANDI, R10,R2,31 //Extracting 5 LSBs of A to find out the value to left rotate by, R11 contains the val
  when x"00000090" => rd <= "001010" & "01010" & "00000" & "00000" & "00000" & "000101";  --BEQ R10, R0, 5 //Skips SHL because R10 is 0
  when x"00000094" => rd <= "000001" & "00000" & "01011" & "00000" & "00000" & "000000";  --ADDI R11,R0,0 //Store 0 for our counter
  when x"00000098" => rd <= "000101" & "00110" & "00110" & "00000" & "00000" & "000001";  --SHL R6,R6,1
  when x"0000009C" => rd <= "000001" & "01011" & "01011" & "00000" & "00000" & "000001";  --ADDI R11, R11, 1 //increment R11
  when x"000000A0" => rd <= "001010" & "01010" & "01011" & "00000" & "00000" & "000001";  --BEQ, R10, R11, 1
  when x"000000A4" => rd <= "001100" & "00000" & "00000" & "00000" & "00000" & "100110";  --JUMP 38 //after the halt
  when x"000000A8" => rd <= "000001" & "00000" & "01100" & "00000" & "00000" & "100000";  --ADDI R12, R0, 32 //R12 = 32
  when x"000000AC" => rd <= "000000" & "01100" & "01010" & "01100" & "00000" & "000011";  --SUB R12, R12, R10 //R12 = 32 - LSB of A
  when x"000000B0" => rd <= "000001" & "00000" & "01101" & "00000" & "00000" & "000000";  --ADDI R13, R0, 0 //R13 = 0 if we are about to right shift B xor A
  when x"000000B4" => rd <= "001100" & "00000" & "00000" & "00000" & "00000" & "111001";  --***CHANGED BY E****JUMP 57 //after the halt
  when x"000000B8" => rd <= "000000" & "00110" & "01110" & "00011" & "00000" & "000001";  --ADD R3, R6, R14 //Adding the left shifted and right shifted components together.
  when x"000000BC" => rd <= "000111" & "00111" & "01000" & "00000" & "00000" & "000001";  --LB R8, R7, 1 //R8 = S[2xi+1]
  when x"000000C0" => rd <= "000000" & "00011" & "01000" & "00011" & "00000" & "000001";  --ADD, R3, R3, R8 //B = ((B xor A) << A) + S[2xi+1]
  when x"000000C4" => rd <= "001000" & "00111" & "00010" & "00000" & "00011" & "000110";  --***ADDED BY E****SB R2, R7, 198 //This should store Mem[2xi + 198] = R2 = A   ----- After 12 rounds this means Mem[200] thorugh Mem[223] should hold all end of
  when x"000000C8" => rd <= "001000" & "00111" & "00011" & "00000" & "00011" & "000111";  --***ADDED BY E****SB R3, R7, 199 //This should store Mem[2xi + 199] = R3 = B
  when x"000000CC" => rd <= "000001" & "00001" & "00001" & "00000" & "00000" & "000001";  --ADDI, R1, R1, 1 //R1 = i = i + 1
  when x"000000D0" => rd <= "001010" & "00001" & "01001" & "00000" & "00000" & "000001";  --BEQ R1, R9, 1 //should loop back to the specified line above
  when x"000000D4" => rd <= "001100" & "00000" & "00000" & "00000" & "00000" & "001000";  --JUMP 8 //after the halt
  when x"000000D8" => rd <= "001000" & "00000" & "00010" & "00000" & "00000" & "011100";  --SB R2, R0, 28
  when x"000000DC" => rd <= "001000" & "00000" & "00011" & "00000" & "00000" & "011101";  --SB R3, R0, 29
  when x"000000E0" => rd <= "111111" & "00000" & "00000" & "00000" & "00000" & "000000";  --HALT
  when x"000000E4" => rd <= "000001" & "00000" & "10010" & "00000" & "00000" & "000000";  --ADDI R18, R0, 0 //R18 is for tracking how many right shifts have been done
  when x"000000E8" => rd <= "000001" & "00000" & "01111" & "00000" & "00000" & "000000";  --ADDI R15, R0, 0 //R15 is for tracking the result of the right shift --- Reg initialized to 0
  when x"000000EC" => rd <= "000111" & "00000" & "10000" & "00000" & "00010" & "000010";  --LB, R16, R0,130 //R16 = Mem(130) = 2147483648
  when x"000000F0" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --BLT R14, R16, 3
  when x"000000F4" => rd <= "000111" & "00000" & "10001" & "00000" & "00010" & "000001";  --LB R17, R0, 129 //R17 = Mem(129) = 1073741824 //R17 to be added to result
  when x"000000F8" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --SUB R14, R14, R16 //a = a - 2147483648
  when x"000000FC" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --ADD R15, R15, R17 //result = result + 1073741824
  when x"00000100" => rd <= "000111" & "00000" & "10000" & "00000" & "00010" & "000001";  --LB, R16, R0,129 //R16 = Mem(129) = 1073741824
  when x"00000104" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --BLT R14, R16, 3
  when x"00000108" => rd <= "000111" & "00000" & "10001" & "00000" & "00010" & "000000";  --LB R17, R0, 128 //R17 = Mem(128) = 536870912 //R17 to hold the amount to be added to result
  when x"0000010C" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --SUB R14, R14, R16 //a = a - 1073741824
  when x"00000110" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --ADD R15, R15, R17 //result = result + 536870912
  when x"00000114" => rd <= "000111" & "00000" & "10000" & "00000" & "00010" & "000000";  --LB, R16, R0,128 //R16 = Mem(128) = 536870912
  when x"00000118" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --BLT R14, R16, 3        
  when x"0000011C" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "111111";  --LB R17, R0, 127 //R17 = Mem(127) = 268435456 //R17 to hold the amount to be added to result
  when x"00000120" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --SUB R14, R14, R16 //a = a - 536870912         
  when x"00000124" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --ADD R15, R15, R17 //result = result + 268435456
  when x"00000128" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "111111";  --LB, R16, R0,127 //R16 = Mem(127) = 268435456
  when x"0000012C" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --BLT R14, R16, 3
  when x"00000130" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "111110";  --LB R17, R0, 126 //R17 = Mem(126) = 134217728 //R17 to hold the amount to be added to result
  when x"00000134" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --SUB R14, R14, R16 //a = a - 268435456
  when x"00000138" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --ADD R15, R15, R17 //result = result + 134217728
  when x"0000013C" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "111110";  --LB, R16, R0,126 //R16 = Mem(126) = 134217728
  when x"00000140" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --BLT R14, R16, 3
  when x"00000144" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "111101";  --LB R17, R0, 125 //R17 = Mem(125) = 67108864 //R17 to hold the amount to be added to result
  when x"00000148" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --SUB R14, R14, R16 //a = a - 134217728
  when x"0000014C" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --ADD R15, R15, R17 //result = result + 67108864
  when x"00000150" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "111101";  --LB, R16, R0,125 //R16 = Mem(125) = 67108864
  when x"00000154" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --BLT R14, R16, 3
  when x"00000158" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "111100";  --LB R17, R0, 124 //R17 = Mem(124) = 33554432 //R17 to hold the amount to be added to result
  when x"0000015C" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --SUB R14, R14, R16 //a = a - 67108864
  when x"00000160" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --ADD R15, R15, R17 //result = result + 33554432
  when x"00000164" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "111100";  --LB, R16, R0,124 //R16 = Mem(124) = 33554432
  when x"00000168" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --BLT R14, R16, 3
  when x"0000016C" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "111011";  --LB R17, R0, 123 //R17 = Mem(123) = 16777216 //R17 to hold the amount to be added to result
  when x"00000170" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --SUB R14, R14, R16 //a = a - 33554432
  when x"00000174" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --ADD R15, R15, R17 //result = result + 16777216
  when x"00000178" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "111011";  --LB, R16, R0,123 //R16 = Mem(123) = 16777216
  when x"0000017C" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --BLT R14, R16, 3
  when x"00000180" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "111010";  --LB R17, R0, 122 //R17 = Mem(122) = 8388608 //R17 to hold the amount to be added to result
  when x"00000184" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --SUB R14, R14, R16 //a = a - 16777216
  when x"00000188" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --ADD R15, R15, R17 //result = result + 8388608
  when x"0000018C" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "111010";  --LB, R16, R0,122 //R16 = Mem(122) = 8388608
  when x"00000190" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --BLT R14, R16, 3
  when x"00000194" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "111001";  --LB R17, R0, 121 //R17 = Mem(121) = 4194304 //R17 to hold the amount to be added to result
  when x"00000198" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --SUB R14, R14, R16 //a = a - 8388608
  when x"0000019C" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --ADD R15, R15, R17 //result = result + 4194304
  when x"000001A0" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "111001";  --LB, R16, R0,121 //R16 = Mem(121) = 4194304
  when x"000001A4" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --BLT R14, R16, 3
  when x"000001A8" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "111000";  --LB R17, R0, 120 //R17 = Mem(120) =  2097152 //R17 to hold the amount to be added to result
  when x"000001AC" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --SUB R14, R14, R16 //a = a - 4194304
  when x"000001B0" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --ADD R15, R15, R17 //result = result +  2097152
  when x"000001B4" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "111000";  --LB, R16, R0,120 //R16 = Mem(120) = 2097152
  when x"000001B8" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --BLT R14, R16, 3
  when x"000001BC" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "110111";  --LB R17, R0, 119 //R17 = Mem(119) = 1048576 //R17 to hold the amount to be added to result
  when x"000001C0" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --SUB R14, R14, R16 //a = a - 2097152
  when x"000001C4" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --ADD R15, R15, R17 //result = result + 1048576
  when x"000001C8" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "110111";  --LB, R16, R0,119 //R16 = Mem(119) = 1048576
  when x"000001CC" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --BLT R14, R16, 3
  when x"000001D0" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "110110";  --LB R17, R0, 118 //R17 = Mem(118) =  524288 //R17 to hold the amount to be added to result
  when x"000001D4" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --SUB R14, R14, R16 //a = a - 1048576
  when x"000001D8" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --ADD R15, R15, R17 //result = result +  524288
  when x"000001DC" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "110110";  --LB, R16, R0,118 //R16 = Mem(118) = 524288
  when x"000001E0" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --BLT R14, R16, 3
  when x"000001E4" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "110101";  --LB R17, R0, 117 //R17 = Mem(117) = 262144 //R17 to hold the amount to be added to result
  when x"000001E8" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --SUB R14, R14, R16 //a = a - 524288
  when x"000001EC" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --ADD R15, R15, R17 //result = result + 262144
  when x"000001F0" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "110101";  --LB, R16, R0,117 //R16 = Mem(117) = 262144
  when x"000001F4" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --BLT R14, R16, 3
  when x"000001F8" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "110100";  --LB R17, R0, 116 //R17 = Mem(116) = 131072 //R17 to hold the amount to be added to result
  when x"000001FC" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --SUB R14, R14, R16 //a = a - 262144
  when x"00000200" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --ADD R15, R15, R17 //result = result + 131072
  when x"00000204" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "110100";  --LB, R16, R0,116 //R16 = Mem(116) = 131072
  when x"00000208" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --BLT R14, R16, 3
  when x"0000020C" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "110011";  --LB R17, R0, 115 //R17 = Mem(115) = 65536 //R17 to hold the amount to be added to result
  when x"00000210" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --SUB R14, R14, R16 //a = a - 131072
  when x"00000214" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --ADD R15, R15, R17 //result = result + 65536
  when x"00000218" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "110011";  --LB, R16, R0,115 //R16 = Mem(115) = 65536
  when x"0000021C" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --BLT R14, R16, 3
  when x"00000220" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "110010";  --LB R17, R0, 114 //R17 = Mem(114) = 32768 //R17 to hold the amount to be added to result
  when x"00000224" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --SUB R14, R14, R16 //a = a - 65536
  when x"00000228" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --ADD R15, R15, R17 //result = result + 32768
  when x"0000022C" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "110010";  --LB, R16, R0,114 //R16 = Mem(114) = 32768
  when x"00000230" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --BLT R14, R16, 3
  when x"00000234" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "110001";  --LB R17, R0, 113 //R17 = Mem(113) = 16384//R17 to hold the amount to be added to result
  when x"00000238" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --SUB R14, R14, R16 //a = a - 32768
  when x"0000023C" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --ADD R15, R15, R17 //result = result + 16384
  when x"00000240" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "110001";  --LB, R16, R0,113 //R16 = Mem(113) = 16384
  when x"00000244" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --BLT R14, R16, 3
  when x"00000248" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "110000";  --LB R17, R0, 112 //R17 = Mem(112) = 8192 //R17 to hold the amount to be added to result
  when x"0000024C" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --SUB R14, R14, R16 //a = a - 16384
  when x"00000250" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --ADD R15, R15, R17 //result = result + 8192
  when x"00000254" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "110000";  --LB, R16, R0,112 //R16 = Mem(112) = 8192
  when x"00000258" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --BLT R14, R16, 3
  when x"0000025C" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "101111";  --LB R17, R0, 111 //R17 = Mem(111) = 4096 //R17 to hold the amount to be added to result
  when x"00000260" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --SUB R14, R14, R16 //a = a - 8192
  when x"00000264" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --ADD R15, R15, R17 //result = result + 4096
  when x"00000268" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "101111";  --LB, R16, R0,111 //R16 = Mem(111) = 4096
  when x"0000026C" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --BLT R14, R16, 3
  when x"00000270" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "101110";  --LB R17, R0, 110 //R17 = Mem(110) = 2048 //R17 to hold the amount to be added to result
  when x"00000274" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --SUB R14, R14, R16 //a = a - 4096
  when x"00000278" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --ADD R15, R15, R17 //result = result + 2048
  when x"0000027C" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "101110";  --LB, R16, R0,110 //R16 = Mem(110) = 2048
  when x"00000280" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --BLT R14, R16, 3
  when x"00000284" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "101101";  --LB R17, R0, 109 //R17 = Mem(109) = 1024 //R17 to hold the amount to be added to result
  when x"00000288" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --SUB R14, R14, R16 //a = a - 2048
  when x"0000028C" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --ADD R15, R15, R17 //result = result + 1024
  when x"00000290" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "101101";  --LB, R16, R0,109 //R16 = Mem(109) = 1024
  when x"00000294" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --BLT R14, R16, 3
  when x"00000298" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "101100";  --LB R17, R0, 108 //R17 = Mem(108) = 512 //R17 to hold the amount to be added to result
  when x"0000029C" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --SUB R14, R14, R16 //a = a - 1024
  when x"000002A0" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --ADD R15, R15, R17 //result = result + 512
  when x"000002A4" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "101100";  --LB, R16, R0,108 //R16 = Mem(108) = 512
  when x"000002A8" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --BLT R14, R16, 3
  when x"000002AC" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "101011";  --LB R17, R0, 107 //R17 = Mem(107) = 256 //R17 to hold the amount to be added to result
  when x"000002B0" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --SUB R14, R14, R16 //a = a - 512
  when x"000002B4" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --ADD R15, R15, R17 //result = result + 256
  when x"000002B8" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "101011";  --LB, R16, R0,107 //R16 = Mem(107) = 256
  when x"000002BC" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --BLT R14, R16, 3
  when x"000002C0" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "101010";  --LB R17, R0, 106 //R17 = Mem(106) = 128 //R17 to hold the amount to be added to result
  when x"000002C4" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --SUB R14, R14, R16 //a = a - 256
  when x"000002C8" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --ADD R15, R15, R17 //result = result + 128
  when x"000002CC" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "101010";  --LB, R16, R0,106 //R16 = Mem(106) = 128
  when x"000002D0" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --BLT R14, R16, 3
  when x"000002D4" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "101001";  --LB R17, R0, 105 //R17 = Mem(105) = 64 //R17 to hold the amount to be added to result
  when x"000002D8" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --SUB R14, R14, R16 //a = a - 128
  when x"000002DC" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --ADD R15, R15, R17 //result = result + 64
  when x"000002E0" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "101001";  --LB, R16, R0,105 //R16 = Mem(105) = 64
  when x"000002E4" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --BLT R14, R16, 3
  when x"000002E8" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "101000";  --LB R17, R0, 104 //R17 = Mem(104) = 32 //R17 to hold the amount to be added to result
  when x"000002EC" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --SUB R14, R14, R16 //a = a - 64
  when x"000002F0" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --ADD R15, R15, R17 //result = result + 32
  when x"000002F4" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "101000";  --LB, R16, R0,104 //R16 = Mem(104) = 32
  when x"000002F8" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --BLT R14, R16, 3
  when x"000002FC" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "100111";  --LB R17, R0, 103 //R17 = Mem(103) = 16 //R17 to hold the amount to be added to result
  when x"00000300" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --SUB R14, R14, R16 //a = a - 32
  when x"00000304" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --ADD R15, R15, R17 //result = result + 16
  when x"00000308" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "100111";  --LB, R16, R0,103 //R16 = Mem(103) = 16
  when x"0000030C" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --BLT R14, R16, 3
  when x"00000310" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "100110";  --LB R17, R0, 102 //R17 = Mem(102) = 8 //R17 to hold the amount to be added to result
  when x"00000314" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --SUB R14, R14, R16 //a = a - 16
  when x"00000318" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --ADD R15, R15, R17 //result = result + 8
  when x"0000031C" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "100110";  --LB, R16, R0,102 //R16 = Mem(102) = 8
  when x"00000320" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --BLT R14, R16, 3
  when x"00000324" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "100101";  --LB R17, R0, 101 //R17 = Mem(101) = 4 //R17 to hold the amount to be added to result
  when x"00000328" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --SUB R14, R14, R16 //a = a - 8
  when x"0000032C" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --ADD R15, R15, R17 //result = result + 4
  when x"00000330" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "100101";  --LB, R16, R0,101 //R16 = Mem(101) = 4
  when x"00000334" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --BLT R14, R16, 3
  when x"00000338" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "100100";  --LB R17, R0, 100 //R17 = Mem(100) = 2 //R17 to hold the amount to be added to result
  when x"0000033C" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --SUB R14, R14, R16 //a = a - 4
  when x"00000340" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --ADD R15, R15, R17 //result = result + 2
  when x"00000344" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "100100";  --LB, R16, R0,100 //R16 = Mem(100) = 2
  when x"00000348" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --BLT R14, R16, 3
  when x"0000034C" => rd <= "000001" & "00000" & "10001" & "00000" & "00000" & "000001";  --ADDI R17, R0, 1 //R17 stores the amount to be added to result
  when x"00000350" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --SUB R14, R14, R16 //a = a - 2
  when x"00000354" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --ADD R15, R15, R17 //result = result + 1
  when x"00000358" => rd <= "000001" & "01111" & "01110" & "00000" & "00000" & "000000";  --ADDI R14, R15, 0 //Store the newly shifted by one value before the next iteration of the loop
  when x"0000035C" => rd <= "000001" & "10010" & "10010" & "00000" & "00000" & "000001";  --ADDI R18, R18, 1 //R18 increments after each single bit right rotate
  when x"00000360" => rd <= "001010" & "01100" & "10010" & "00000" & "00000" & "000001";  --BEQ R18, R12, 1 //If we've shifted right enough times, skip the jump
  when x"00000364" => rd <= "001100" & "00000" & "00000" & "00000" & "00000" & "111010";  --***CHANGED BY E****JUMP 58 //should jump to after the initialization period of the right shift
  when x"00000368" => rd <= "001010" & "00000" & "01101" & "00000" & "00000" & "000001";  --BEQ R13, R0, //branch back to after the B xor A left rotate
  when x"0000036C" => rd <= "001100" & "00000" & "00000" & "00000" & "00000" & "011001";  --JUMP 25 //Jump back to after the A xor B left rotate
  when x"00000370" => rd <= "001100" & "00000" & "00000" & "00000" & "00000" & "101110";  --JUMP 46
  when others  => rd <= (others => '0');         
end case;
end process;

end rtl;