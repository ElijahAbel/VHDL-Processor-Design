library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity instructMem is
port (
  instructAddr : in std_logic_vector(31 downto 0); --input instruction from PC
  rd           : out std_logic_vector(31 downto 0) --output instruction to decoder and register file
);
end instructMem;

architecture rtl of instructMem is

-- --OPCODES
-- signal ARITH    : std_logic_vector(5 downto 0) := "000000"; --OPCODE00
-- signal ADDIMM   : std_logic_vector(5 downto 0) := "000001"; --OPCODE01
-- signal SUBIMM   : std_logic_vector(5 downto 0) := "000010"; --OPCODE02
-- signal ANDIMM   : std_logic_vector(5 downto 0) := "000011"; --OPCODE03
-- signal ORIMM    : std_logic_vector(5 downto 0) := "000100"; --OPCODE04
-- signal SHFLFT   : std_logic_vector(5 downto 0) := "000101"; --OPCODE05
-- signal LOAD     : std_logic_vector(5 downto 0) := "000111"; --OPCODE07
-- signal STORE    : std_logic_vector(5 downto 0) := "001000"; --OPCODE08
-- signal BLT      : std_logic_vector(5 downto 0) := "001001"; --OPCODE09
-- signal BEQ      : std_logic_vector(5 downto 0) := "001010"; --OPCODE0A
-- signal BNE      : std_logic_vector(5 downto 0) := "001011"; --OPCODE0B
-- signal JUMP     : std_logic_vector(5 downto 0) := "001100"; --OPCODE0C
-- signal HALT     : std_logic_vector(5 downto 0) := "111111"; --OPCODE3F

-- --FUNCTIONS
-- signal ADDREG   : std_logic_vector(5 downto 0) := "000001"; --FUNC1
-- signal SUBREG   : std_logic_vector(5 downto 0) := "000011"; --FUNC3
-- signal ANDREG   : std_logic_vector(5 downto 0) := "000101"; --FUNC5
-- signal ORREG    : std_logic_vector(5 downto 0) := "000111"; --FUNC7
-- signal NORREG   : std_logic_vector(5 downto 0) := "001001"; --FUNC9

begin

instruct : process (instructAddr)
begin
case instructAddr(31 downto 0) is
                            -- OPCODE&   RS    &  RT     &  RD     &  SHAMT  & FUNCT (R-TYPE)
				            -- OPCODE&   RS    &  RT     & Address/Immediate         (I-TYPE)
				            -- OPCODE&   Address (26-bits)                           (J-TYPE)
  when x"00000000" => rd <= "000000" & "00000" & "00000" & "00000" & "00000" & "000011";  --0   SUB R0, R0, R0     ----- initialize R0 to be 0
  when x"00000004" => rd <= "000000" & "00100" & "00100" & "00100" & "00000" & "000011";  --1   SUB R4, R4, R4
  when x"00000008" => rd <= "000000" & "11011" & "11011" & "11011" & "00000" & "000011";  --2   SUB R27, R27, R27
  when x"0000000C" => rd <= "000001" & "00000" & "11001" & "00000" & "00000" & "000100";  --3   ADDI R25 R0 4
  when x"00000010" => rd <= "000001" & "00000" & "01000" & "00000" & "00001" & "111111";  --4   ADDI R8, R0, 127
  when x"00000014" => rd <= "000000" & "11000" & "11000" & "11000" & "00000" & "000011";  --5   SUB R24, R24, R24
  when x"00000018" => rd <= "000000" & "11010" & "11010" & "11010" & "00000" & "000011";  --6   SUB R26, R26, R26
  when x"0000001C" => rd <= "001011" & "11000" & "11001" & "00000" & "00000" & "000011";  --7   BNE R24, R25, 4    --**BPa   
  when x"00000020" => rd <= "000001" & "11010" & "11010" & "00000" & "00000" & "000001";  --8   ADDI R26, R26, 1
  when x"00000024" => rd <= "001010" & "11001" & "11010" & "00000" & "00000" & "001101";  --9   BEQ R26, R25, 13
  when x"00000028" => rd <= "000000" & "11000" & "11000" & "11000" & "00000" & "000011";  --10  SUB R24, R24, R24
  when x"0000002C" => rd <= "000111" & "11010" & "00111" & "00000" & "00000" & "110010";  --11  LW  R7,50(R26) 
  when x"00000030" => rd <= "000000" & "00111" & "01000" & "01001" & "00000" & "000101";  --12  AND R9 R8 R7
  when x"00000034" => rd <= "000101" & "00011" & "00011" & "00000" & "00000" & "001000";  --13  SHL R3, R3, 8
  when x"00000038" => rd <= "000000" & "00011" & "01001" & "00011" & "00000" & "000001";  --14  ADD R3 R9 R3
  when x"0000003C" => rd <= "001000" & "11000" & "00011" & "00000" & "00000" & "110111";  --15  SW  R3,55(R26)
  when x"00000040" => rd <= "000101" & "00111" & "00110" & "00000" & "00000" & "001000";  --16  SHL R6,R7, 8  
  when x"00000044" => rd <= "000001" & "00111" & "01110" & "00000" & "00000" & "000000";  --17  ADDI R14, R7, 0 
  when x"00000048" => rd <= "000001" & "00000" & "10011" & "00000" & "00000" & "011000";  --18  ADDI R19, R0, 24 
  when x"0000004C" => rd <= "001100" & "00000" & "00000" & "00000" & "00001" & "111111";  --19  JMP  127
  when x"00000050" => rd <= "000000" & "00110" & "01111" & "00111" & "00000" & "000001";  --20  ADD R7, R6, R15 
  when x"00000054" => rd <= "000001" & "11000" & "11000" & "00000" & "00000" & "000001";  --21  ADDI R24, R24, 1  
  when x"00000058" => rd <= "001100" & "00000" & "00000" & "00000" & "00000" & "000111";  --22  JMP   7
  when x"0000005C" => rd <= "000001" & "00000" & "01010" & "10110" & "11111" & "100001";  --23  ADDI R10, R0, hex(B7E1)      -- assign Pw to R10, Qw to R11
  when x"00000060" => rd <= "000101" & "01010" & "01010" & "00000" & "00000" & "010000";  --24  SHL R10, R10, 16
  when x"00000064" => rd <= "000001" & "01010" & "01010" & "01010" & "00101" & "100011";  --25  ADDI R10, R10, hex(5163)
  when x"00000068" => rd <= "000001" & "00000" & "01011" & "10011" & "11000" & "110111";  --26  ADDI R11, R0, hex(9E37)
  when x"0000006C" => rd <= "000101" & "01011" & "01011" & "00000" & "00000" & "010000";  --27  SHL R11, R11, 16
  when x"00000070" => rd <= "000001" & "01011" & "01011" & "01111" & "00110" & "111001";  --28  ADDI R11, R11, hex(79B9)
  when x"00000074" => rd <= "001000" & "00000" & "01010" & "00000" & "00000" & "111100";  --29  SW  R10, 60(R0)
  when x"00000078" => rd <= "000000" & "01010" & "01011" & "01010" & "00000" & "000001";  --30  ADD R10, R11, R10
  when x"0000007C" => rd <= "001000" & "00000" & "01010" & "00000" & "00000" & "111101";  --31  SW  R10, 61(R0)
  when x"00000080" => rd <= "000000" & "01010" & "01011" & "01010" & "00000" & "000001";  --32  ADD R10, R11, R10
  when x"00000084" => rd <= "001000" & "00000" & "01010" & "00000" & "00000" & "111110";  --33  SW  R10, 62(R0)
  when x"00000088" => rd <= "000000" & "01010" & "01011" & "01010" & "00000" & "000001";  --34  ADD R10, R11, R10
  when x"0000008C" => rd <= "001000" & "00000" & "01010" & "00000" & "00000" & "111111";  --35  SW  R10, 63(R0)
  when x"00000090" => rd <= "000000" & "01010" & "01011" & "01010" & "00000" & "000001";  --36  ADD R10, R11, R10
  when x"00000094" => rd <= "001000" & "00000" & "01010" & "00000" & "00001" & "000000";  --37  SW  R10, 64(R0)
  when x"00000098" => rd <= "000000" & "01010" & "01011" & "01010" & "00000" & "000001";  --38  ADD R10, R11, R10
  when x"0000009C" => rd <= "001000" & "00000" & "01010" & "00000" & "00001" & "000001";  --39  SW  R10, 65(R0)
  when x"000000A0" => rd <= "000000" & "01010" & "01011" & "01010" & "00000" & "000001";  --40  ADD R10, R11, R10
  when x"000000A4" => rd <= "001000" & "00000" & "01010" & "00000" & "00001" & "000010";  --41  SW  R10, 66(R0)
  when x"000000A8" => rd <= "000000" & "01010" & "01011" & "01010" & "00000" & "000001";  --42  ADD R10, R11, R10
  when x"000000AC" => rd <= "001000" & "00000" & "01010" & "00000" & "00001" & "000011";  --43  SW  R10, 67(R0)
  when x"000000B0" => rd <= "000000" & "01010" & "01011" & "01010" & "00000" & "000001";  --44  ADD R10, R11, R10
  when x"000000B4" => rd <= "001000" & "00000" & "01010" & "00000" & "00001" & "000100";  --45  SW  R10, 68(R0)
  when x"000000B8" => rd <= "000000" & "01010" & "01011" & "01010" & "00000" & "000001";  --46  ADD R10, R11, R10
  when x"000000BC" => rd <= "001000" & "00000" & "01010" & "00000" & "00001" & "000101";  --47  SW  R10, 69(R0)
  when x"000000C0" => rd <= "000000" & "01010" & "01011" & "01010" & "00000" & "000001";  --48  ADD R10, R11, R10
  when x"000000C4" => rd <= "001000" & "00000" & "01010" & "00000" & "00001" & "000110";  --49  SW  R10, 70(R0)em[223] should hold all end of
  when x"000000C8" => rd <= "000000" & "01010" & "01011" & "01010" & "00000" & "000001";  --50  ADD R10, R11, R10
  when x"000000CC" => rd <= "001000" & "00000" & "01010" & "00000" & "00001" & "000111";  --51  SW  R10, 71(R0)
  when x"000000D0" => rd <= "000000" & "01010" & "01011" & "01010" & "00000" & "000001";  --52  ADD R10, R11, R10
  when x"000000D4" => rd <= "001000" & "00000" & "01010" & "00000" & "00001" & "001000";  --53  SW  R10, 72(R0)
  when x"000000D8" => rd <= "000000" & "01010" & "01011" & "01010" & "00000" & "000001";  --54  ADD R10, R11, R10
  when x"000000DC" => rd <= "001000" & "00000" & "01010" & "00000" & "00001" & "001001";  --55  SW  R10, 73(R0)
  when x"000000E0" => rd <= "000000" & "01010" & "01011" & "01010" & "00000" & "000001";  --56  ADD R10, R11, R10
  when x"000000E4" => rd <= "001000" & "00000" & "01010" & "00000" & "00001" & "001010";  --57  SW  R10, 74(R0)
  when x"000000E8" => rd <= "000000" & "01010" & "01011" & "01010" & "00000" & "000001";  --58  ADD R10, R11, R10
  when x"000000EC" => rd <= "001000" & "00000" & "01010" & "00000" & "00001" & "001011";  --59  SW  R10, 75(R0)
  when x"000000F0" => rd <= "000000" & "01010" & "01011" & "01010" & "00000" & "000001";  --60  ADD R10, R11, R10
  when x"000000F4" => rd <= "001000" & "00000" & "01010" & "00000" & "00001" & "001100";  --61  SW  R10, 76(R0)
  when x"000000F8" => rd <= "000000" & "01010" & "01011" & "01010" & "00000" & "000001";  --62  ADD R10, R11, R10
  when x"000000FC" => rd <= "001000" & "00000" & "01010" & "00000" & "00001" & "001101";  --63  SW  R10, 77(R0)
  when x"00000100" => rd <= "000000" & "01010" & "01011" & "01010" & "00000" & "000001";  --64  ADD R10, R11, R10
  when x"00000104" => rd <= "001000" & "00000" & "01010" & "00000" & "00001" & "001110";  --65  SW  R10, 78(R0)
  when x"00000108" => rd <= "000000" & "01010" & "01011" & "01010" & "00000" & "000001";  --66  ADD R10, R11, R10
  when x"0000010C" => rd <= "001000" & "00000" & "01010" & "00000" & "00001" & "001111";  --67  SW  R10, 79(R0)
  when x"00000110" => rd <= "000000" & "01010" & "01011" & "01010" & "00000" & "000001";  --68  ADD R10, R11, R10
  when x"00000114" => rd <= "001000" & "00000" & "01010" & "00000" & "00001" & "010000";  --69  SW  R10, 80(R0)
  when x"00000118" => rd <= "000000" & "01010" & "01011" & "01010" & "00000" & "000001";  --70  ADD R10, R11, R10
  when x"0000011C" => rd <= "001000" & "00000" & "01010" & "00000" & "00001" & "010001";  --71  SW  R10, 81(R0)
  when x"00000120" => rd <= "000000" & "01010" & "01011" & "01010" & "00000" & "000001";  --72  ADD R10, R11, R10
  when x"00000124" => rd <= "001000" & "00000" & "01010" & "00000" & "00001" & "010010";  --73  SW  R10, 82(R0)
  when x"00000128" => rd <= "000000" & "01010" & "01011" & "01010" & "00000" & "000001";  --74  ADD R10, R11, R10
  when x"0000012C" => rd <= "001000" & "00000" & "01010" & "00000" & "00001" & "010011";  --75  SW  R10, 83(R0)
  when x"00000130" => rd <= "000000" & "01010" & "01011" & "01010" & "00000" & "000001";  --76  ADD R10, R11, R10
  when x"00000134" => rd <= "001000" & "00000" & "01010" & "00000" & "00001" & "010100";  --77  SW  R10, 84(R0)
  when x"00000138" => rd <= "000000" & "01010" & "01011" & "01010" & "00000" & "000001";  --78  ADD R10, R11, R10
  when x"0000013C" => rd <= "001000" & "00000" & "01010" & "00000" & "00001" & "010101";  --79  SW  R10, 85(R0)
  when x"00000140" => rd <= "000000" & "11011" & "11011" & "11011" & "00000" & "000011";  --80  SUB R27, R27, R27
  when x"00000144" => rd <= "000001" & "00000" & "00100" & "00000" & "00000" & "011010";  --81  ADDI R4, R0, 26   -- R14 = t = 26
  when x"00000148" => rd <= "000001" & "00000" & "00101" & "00000" & "00000" & "000100";  --82  ADDI R5, R0, 4    -- R15 = c = 4
  when x"0000014C" => rd <= "000000" & "00001" & "00001" & "00001" & "00000" & "000011";  --83  SUB R1, R1, R1     -- clear R1 and R2 to be 0
  when x"00000150" => rd <= "000000" & "00010" & "00010" & "00010" & "00000" & "000011";  --84  SUB R2, R2, R2     -- For A and B ( initial values are 0)
  when x"00000154" => rd <= "000000" & "01010" & "01010" & "01010" & "00000" & "000011";  --85  SUB R10, R10, R10  --  i = 0
  when x"00000158" => rd <= "000000" & "01011" & "01011" & "01011" & "00000" & "000011";  --86  SUB R11, R11, R11  --  j = 0
  when x"0000015C" => rd <= "000001" & "11110" & "11110" & "00000" & "00001" & "001110";  --87  ADDI R30, R30, 78
  when x"00000160" => rd <= "000000" & "11111" & "11111" & "11111" & "00000" & "000011";  --88  SUB R31, R31, R31  --  if R31 == 78, we stop
  when x"00000164" => rd <= "001011" & "11110" & "11111" & "00000" & "00000" & "000011";  --89  BNE R30, R31, 3    --  the start of the loop
  when x"00000168" => rd <= "001000" & "00000" & "00001" & "00000" & "00001" & "011010";  --90  SW  R1, 90(R0)       -- Assuming A will be stored to Mem[90]
  when x"0000016C" => rd <= "001000" & "00000" & "00010" & "00000" & "00001" & "011011";  --91  SW  R2, 91(R0)       -- Assuming B will be stored to Mem[91]
  when x"00000170" => rd <= "111111" & "00000" & "00000" & "00000" & "00000" & "000000";  --92  HLT
  when x"00000174" => rd <= "000001" & "11111" & "11111" & "00000" & "00000" & "000001";  --93  ADDI R31,R31,1
  when x"00000178" => rd <= "000111" & "01010" & "01100" & "00000" & "00000" & "111100";  --94  LW  R12, 60(R10)
  when x"0000017C" => rd <= "000000" & "01100" & "00001" & "01100" & "00000" & "000001";  --95  ADD R12, R1, R12
  when x"00000180" => rd <= "000000" & "01100" & "00010" & "01100" & "00000" & "000001";  --96  ADD R12, R2, R12
  when x"00000184" => rd <= "000101" & "01100" & "00110" & "00000" & "00000" & "000011";  --97  SHL R6,R12, 3     ---- storing the left shift part to R6
  when x"00000188" => rd <= "000001" & "01100" & "01110" & "00000" & "00000" & "000000";  --98  ADDI R14, R12, 0  ---- storing the original value to R14
  when x"0000018C" => rd <= "000001" & "00000" & "10011" & "00000" & "00000" & "011101";  --99  ADDI R19, R0, 29  ----- R19 is bits for right shift
  when x"00000190" => rd <= "001100" & "00000" & "00000" & "00000" & "00001" & "111111";  --100 JMP 127 (RIght shift)
  when x"00000194" => rd <= "000000" & "00110" & "01111" & "01100" & "00000" & "000001";  --101 ADD R12, R6, R15   ---- back point   (BP1)
  when x"00000198" => rd <= "001000" & "01010" & "01100" & "00000" & "00000" & "111100";  --102 SW  R12, 60(R10)
  when x"0000019C" => rd <= "000000" & "01100" & "00000" & "00001" & "00000" & "000001";  --103 ADD R1, R12, R0
  when x"000001A0" => rd <= "000111" & "01011" & "01101" & "00000" & "00000" & "110111";  --104 LW  R13, 55(R11)       --
  when x"000001A4" => rd <= "000000" & "00001" & "00010" & "00010" & "00000" & "000001";  --105 ADD R2, R1, R2        --R2 stores A + B, which is also the times we need to shift
  when x"000001A8" => rd <= "000000" & "00010" & "01101" & "01101" & "00000" & "000001";  --106 ADD R13, R2, R13
  when x"000001AC" => rd <= "000001" & "01101" & "01110" & "00000" & "00000" & "000000";  --107 ADDI R14, R13, 0
  when x"000001B0" => rd <= "000001" & "00000" & "01000" & "00000" & "00000" & "011111";  --108 ADDI R8, R0, 32
  when x"000001B4" => rd <= "000000" & "00010" & "01000" & "00110" & "00000" & "000101";  --109 AND  R6, R2, R8    ---   R6 : bits to left shift
  when x"000001B8" => rd <= "000001" & "00000" & "10011" & "00000" & "00000" & "100000";  --110 ADDI R19, R0, 32
  when x"000001BC" => rd <= "000000" & "10011" & "00110" & "10011" & "00000" & "000011";  --111 SUB  R19, R19, R6  ----  R19 : bits to righ shift
  when x"000001C0" => rd <= "001010" & "00110" & "00000" & "00000" & "00000" & "000011";  --112 BEQ R6, R0, 3
  when x"000001C4" => rd <= "000101" & "01101" & "01101" & "00000" & "00000" & "000001";  --113 SHL R13, R13, 1
  when x"000001C8" => rd <= "000010" & "00110" & "00110" & "00000" & "00000" & "000001";  --114 SUBI R6, R6, 1
  when x"000001CC" => rd <= "001100" & "00000" & "00000" & "00000" & "00001" & "110000";  --115 JMP 112######
  when x"000001D0" => rd <= "001100" & "00000" & "00000" & "00000" & "00001" & "111111";  --116 JMP 127  (RIGHT SHIFT)
  when x"000001D4" => rd <= "000000" & "01111" & "01101" & "01101" & "00000" & "000001";  --117 ADD R13, R13, R15    ------   BP2 
  when x"000001D8" => rd <= "000000" & "01101" & "00000" & "00010" & "00000" & "000001";  --118 ADD R2, R13, R0
  when x"000001DC" => rd <= "001000" & "01011" & "00010" & "00000" & "00000" & "110111";  --119 SW  R2, 55(R11)
  when x"000001E0" => rd <= "000001" & "01010" & "01010" & "00000" & "00000" & "000001";  --120 ADDI R10, R10, 1
  when x"000001E4" => rd <= "000001" & "01011" & "01011" & "00000" & "00000" & "000001";  --121 ADDI R11, R11, 1
  when x"000001E8" => rd <= "001011" & "01010" & "00100" & "00000" & "00000" & "000001";  --122 BNE R10, R4, 1      -- i==t and j==c can't be true simutaneously
  when x"000001EC" => rd <= "000000" & "01010" & "01010" & "01010" & "00000" & "000011";  --123 SUB R10, R10, R10
  when x"000001F0" => rd <= "001011" & "01011" & "00101" & "00000" & "00000" & "000001";  --124 BNE R11, R5, 1
  when x"000001F4" => rd <= "000000" & "01011" & "01011" & "01011" & "00000" & "000011";  --125 SUB R11, R11, R11    --  reset R11 = i = 0
  when x"000001F8" => rd <= "001100" & "00000" & "00000" & "00000" & "00001" & "011001";  --126 JMP 89
  when x"000001FC" => rd <= "000001" & "00000" & "10010" & "00000" & "00000" & "000000";  --127 ***RIGHT SHIFT*** --ADDI R18, R0, 0
  when x"00000200" => rd <= "000001" & "00000" & "01111" & "00000" & "00000" & "000000";  --128 *** BP0 *** --ADDI R15, R0, 0 
  when x"00000204" => rd <= "000111" & "00000" & "10000" & "00000" & "00010" & "000010";  --129 LB, R16, R0,130
  when x"00000208" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --130 BLT R14, R16, 3
  when x"0000020C" => rd <= "000111" & "00000" & "10001" & "00000" & "00010" & "000001";  --131 LB R17, R0, 129 
  when x"00000210" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --132 SUB R14, R14, R16
  when x"00000214" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --133 ADD R15, R15, R17 //result = result + 1073741824
  when x"00000218" => rd <= "000111" & "00000" & "10000" & "00000" & "00010" & "000001";  --134 LB, R16, R0,129 //R16 = Mem(129) = 1073741824
  when x"0000021C" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --135 BLT R14, R16, 3
  when x"00000220" => rd <= "000111" & "00000" & "10001" & "00000" & "00010" & "000000";  --136 LB R17, R0, 128 //R17 = Mem(128) = 536870912 //R17 to hold the amount to be added to result
  when x"00000224" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --137 SUB R14, R14, R16 //a = a - 1073741824
  when x"00000228" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --138 ADD R15, R15, R17 //result = result + 536870912
  when x"0000022C" => rd <= "000111" & "00000" & "10000" & "00000" & "00010" & "000000";  --139 LB, R16, R0,128 //R16 = Mem(128) = 536870912
  when x"00000230" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --140 BLT R14, R16, 3        
  when x"00000234" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "111111";  --141 LB R17, R0, 127 //R17 = Mem(127) = 268435456 //R17 to hold the amount to be added to result
  when x"00000238" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --142 SUB R14, R14, R16 //a = a - 536870912         
  when x"0000023C" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --143 ADD R15, R15, R17 //result = result + 268435456
  when x"00000240" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "111111";  --144 LB, R16, R0,127 //R16 = Mem(127) = 268435456
  when x"00000244" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --145 BLT R14, R16, 3
  when x"00000248" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "111110";  --146 LB R17, R0, 126 //R17 = Mem(126) = 134217728 //R17 to hold the amount to be added to result
  when x"0000024C" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --147 SUB R14, R14, R16 //a = a - 268435456
  when x"00000250" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --148 ADD R15, R15, R17 //result = result + 134217728
  when x"00000254" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "111110";  --149 LB, R16, R0,126 //R16 = Mem(126) = 134217728
  when x"00000258" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --150 BLT R14, R16, 3
  when x"0000025C" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "111101";  --151 LB R17, R0, 125 //R17 = Mem(125) = 67108864 //R17 to hold the amount to be added to result
  when x"00000260" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --152 SUB R14, R14, R16 //a = a - 134217728
  when x"00000264" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --153 ADD R15, R15, R17 //result = result + 67108864
  when x"00000268" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "111101";  --154 LB, R16, R0,125 //R16 = Mem(125) = 67108864
  when x"0000026C" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --155 BLT R14, R16, 3
  when x"00000270" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "111100";  --156 LB R17, R0, 124 //R17 = Mem(124) = 33554432 //R17 to hold the amount to be added to result
  when x"00000274" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --157 SUB R14, R14, R16 //a = a - 67108864
  when x"00000278" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --158 ADD R15, R15, R17 //result = result + 33554432
  when x"0000027C" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "111100";  --159 LB, R16, R0,124 //R16 = Mem(124) = 33554432
  when x"00000280" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --160 BLT R14, R16, 3
  when x"00000284" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "111011";  --161 LB R17, R0, 123 //R17 = Mem(123) = 16777216 //R17 to hold the amount to be added to result
  when x"00000288" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --162 SUB R14, R14, R16 //a = a - 33554432
  when x"0000028C" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --163 ADD R15, R15, R17 //result = result + 16777216
  when x"00000290" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "111011";  --164 LB, R16, R0,123 //R16 = Mem(123) = 16777216
  when x"00000294" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --165 BLT R14, R16, 3
  when x"00000298" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "111010";  --166 LB R17, R0, 122 //R17 = Mem(122) = 8388608 //R17 to hold the amount to be added to result
  when x"0000029C" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --167 SUB R14, R14, R16 //a = a - 16777216
  when x"000002A0" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --168 ADD R15, R15, R17 //result = result + 8388608
  when x"000002A4" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "111010";  --169 LB, R16, R0,122 //R16 = Mem(122) = 8388608
  when x"000002A8" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --170 BLT R14, R16, 3
  when x"000002AC" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "111001";  --171 LB R17, R0, 121 //R17 = Mem(121) = 4194304 //R17 to hold the amount to be added to result
  when x"000002B0" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --172 SUB R14, R14, R16 //a = a - 8388608
  when x"000002B4" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --173 ADD R15, R15, R17 //result = result + 4194304
  when x"000002B8" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "111001";  --174 LB, R16, R0,121 //R16 = Mem(121) = 4194304
  when x"000002BC" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --175 BLT R14, R16, 3
  when x"000002C0" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "111000";  --176 LB R17, R0, 120 //R17 = Mem(120) =  2097152 //R17 to hold the amount to be added to result
  when x"000002C4" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --177 SUB R14, R14, R16 //a = a - 4194304
  when x"000002C8" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --178 ADD R15, R15, R17 //result = result +  2097152
  when x"000002CC" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "111000";  --179 LB, R16, R0,120 //R16 = Mem(120) = 2097152
  when x"000002D0" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --180 BLT R14, R16, 3
  when x"000002D4" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "110111";  --181 LB R17, R0, 119 //R17 = Mem(119) = 1048576 //R17 to hold the amount to be added to result
  when x"000002D8" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --182 SUB R14, R14, R16 //a = a - 2097152
  when x"000002DC" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --183 ADD R15, R15, R17 //result = result + 1048576
  when x"000002E0" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "110111";  --184 LB, R16, R0,119 //R16 = Mem(119) = 1048576
  when x"000002E4" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --185 BLT R14, R16, 3
  when x"000002E8" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "110110";  --186 LB R17, R0, 118 //R17 = Mem(118) =  524288 //R17 to hold the amount to be added to result
  when x"000002EC" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --187 SUB R14, R14, R16 //a = a - 1048576
  when x"000002F0" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --188 ADD R15, R15, R17 //result = result +  524288
  when x"000002F4" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "110110";  --189 LB, R16, R0,118 //R16 = Mem(118) = 524288
  when x"000002F8" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --190 BLT R14, R16, 3
  when x"000002FC" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "110101";  --191 LB R17, R0, 117 //R17 = Mem(117) = 262144 //R17 to hold the amount to be added to result
  when x"00000300" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --192 SUB R14, R14, R16 //a = a - 524288
  when x"00000304" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --193 ADD R15, R15, R17 //result = result + 262144
  when x"00000308" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "110101";  --194 LB, R16, R0,117 //R16 = Mem(117) = 262144
  when x"0000030C" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --195 BLT R14, R16, 3
  when x"00000310" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "110100";  --196 LB R17, R0, 116 //R17 = Mem(116) = 131072 //R17 to hold the amount to be added to result
  when x"00000314" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --197 SUB R14, R14, R16 //a = a - 262144
  when x"00000318" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --198 ADD R15, R15, R17 //result = result + 131072
  when x"0000031C" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "110100";  --199 LB, R16, R0,116 //R16 = Mem(116) = 131072
  when x"00000320" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --100 BLT R14, R16, 3
  when x"00000324" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "110011";  --201 LB R17, R0, 115 //R17 = Mem(115) = 65536 //R17 to hold the amount to be added to result
  when x"00000328" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --202 SUB R14, R14, R16 //a = a - 131072
  when x"0000032C" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --203 ADD R15, R15, R17 //result = result + 65536
  when x"00000330" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "110011";  --204 LB, R16, R0,115 //R16 = Mem(115) = 65536
  when x"00000334" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --205 BLT R14, R16, 3
  when x"00000338" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "110010";  --206 LB R17, R0, 114 //R17 = Mem(114) = 32768 //R17 to hold the amount to be added to result
  when x"0000033C" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --207 SUB R14, R14, R16 //a = a - 65536
  when x"00000340" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --208 ADD R15, R15, R17 //result = result + 32768
  when x"00000344" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "110010";  --209 LB, R16, R0,114 //R16 = Mem(114) = 32768
  when x"00000348" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --210 BLT R14, R16, 3
  when x"0000034C" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "110001";  --211 LB R17, R0, 113 //R17 = Mem(113) = 16384//R17 to hold the amount to be added to result
  when x"00000350" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --212 SUB R14, R14, R16 //a = a - 32768
  when x"00000354" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --213 ADD R15, R15, R17 //result = result + 16384
  when x"00000358" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "110001";  --214 LB, R16, R0,113 //R16 = Mem(113) = 16384
  when x"0000035C" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --215 BLT R14, R16, 3
  when x"00000360" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "110000";  --216 LB R17, R0, 112 //R17 = Mem(112) = 8192 //R17 to hold the amount to be added to result
  when x"00000364" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --217 SUB R14, R14, R16 //a = a - 16384
  when x"00000368" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --218 ADD R15, R15, R17 //result = result + 8192
  when x"0000036C" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "110000";  --219 LB, R16, R0,112 //R16 = Mem(112) = 8192
  when x"00000370" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --220 BLT R14, R16, 3
  when x"00000374" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "101111";  --221 LB R17, R0, 111 //R17 = Mem(111) = 4096 //R17 to hold the amount to be added to result
  when x"00000378" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --222 SUB R14, R14, R16 //a = a - 8192
  when x"0000037C" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --223 ADD R15, R15, R17 //result = result + 4096
  when x"00000380" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "101111";  --224 LB, R16, R0,111 //R16 = Mem(111) = 4096
  when x"00000384" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --225 BLT R14, R16, 3
  when x"00000388" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "101110";  --226 LB R17, R0, 110 //R17 = Mem(110) = 2048 //R17 to hold the amount to be added to result
  when x"0000038C" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --227 SUB R14, R14, R16 //a = a - 4096
  when x"00000390" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --228 ADD R15, R15, R17 //result = result + 2048
  when x"00000394" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "101110";  --229 LB, R16, R0,110 //R16 = Mem(110) = 2048
  when x"00000398" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --230 BLT R14, R16, 3
  when x"0000039C" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "101101";  --231 LB R17, R0, 109 //R17 = Mem(109) = 1024 //R17 to hold the amount to be added to result
  when x"000003A0" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --232 SUB R14, R14, R16 //a = a - 2048
  when x"000003A4" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --233 ADD R15, R15, R17 //result = result + 1024
  when x"000003A8" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "101101";  --234 LB, R16, R0,109 //R16 = Mem(109) = 1024
  when x"000003AC" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --235 BLT R14, R16, 3
  when x"000003B0" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "101100";  --236 LB R17, R0, 108 //R17 = Mem(108) = 512 //R17 to hold the amount to be added to result
  when x"000003B4" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --237 SUB R14, R14, R16 //a = a - 1024
  when x"000003B8" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --238 ADD R15, R15, R17 //result = result + 512
  when x"000003BC" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "101100";  --239 LB, R16, R0,108 //R16 = Mem(108) = 512
  when x"000003C0" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --240 BLT R14, R16, 3
  when x"000003C4" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "101011";  --241 LB R17, R0, 107 //R17 = Mem(107) = 256 //R17 to hold the amount to be added to result
  when x"000003C8" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --242 SUB R14, R14, R16 //a = a - 512
  when x"000003CC" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --243 ADD R15, R15, R17 //result = result + 256
  when x"000003D0" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "101011";  --244 LB, R16, R0,107 //R16 = Mem(107) = 256
  when x"000003D4" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --245 BLT R14, R16, 3
  when x"000003D8" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "101010";  --246 LB R17, R0, 106 //R17 = Mem(106) = 128 //R17 to hold the amount to be added to result
  when x"000003DC" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --247 SUB R14, R14, R16 //a = a - 256
  when x"000003E0" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --248 ADD R15, R15, R17 //result = result + 128
  when x"000003E4" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "101010";  --249 LB, R16, R0,106 //R16 = Mem(106) = 128
  when x"000003E8" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --250 BLT R14, R16, 3
  when x"000003EC" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "101001";  --251 LB R17, R0, 105 //R17 = Mem(105) = 64 //R17 to hold the amount to be added to result
  when x"000003F0" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --252 SUB R14, R14, R16 //a = a - 128
  when x"000003F4" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --253 ADD R15, R15, R17 //result = result + 64
  when x"000003F8" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "101001";  --254 LB, R16, R0,105 //R16 = Mem(105) = 64
  when x"000003FC" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --255 BLT R14, R16, 3
  when x"00000400" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "101000";  --256 LB R17, R0, 104 //R17 = Mem(104) = 32 //R17 to hold the amount to be added to result
  when x"00000404" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --257 SUB R14, R14, R16 //a = a - 64
  when x"00000408" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --258 ADD R15, R15, R17 //result = result + 32
  when x"0000040C" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "101000";  --259 LB, R16, R0,104 //R16 = Mem(104) = 32
  when x"00000410" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --260 BLT R14, R16, 3
  when x"00000414" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "100111";  --261 LB R17, R0, 103 //R17 = Mem(103) = 16 //R17 to hold the amount to be added to result
  when x"00000418" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --262 SUB R14, R14, R16 //a = a - 32
  when x"0000041C" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --263 ADD R15, R15, R17 //result = result + 16
  when x"00000420" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "100111";  --264 LB, R16, R0,103 //R16 = Mem(103) = 16
  when x"00000424" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --265 BLT R14, R16, 3
  when x"00000428" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "100110";  --266 LB R17, R0, 102 //R17 = Mem(102) = 8 //R17 to hold the amount to be added to result
  when x"0000042C" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --267 SUB R14, R14, R16 //a = a - 16
  when x"00000430" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --268 ADD R15, R15, R17 //result = result + 8
  when x"00000434" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "100110";  --269 LB, R16, R0,102 //R16 = Mem(102) = 8
  when x"00000438" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --270 BLT R14, R16, 3
  when x"0000043C" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "100101";  --271 LB R17, R0, 101 //R17 = Mem(101) = 4 //R17 to hold the amount to be added to result
  when x"00000440" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --272 SUB R14, R14, R16 //a = a - 8
  when x"00000444" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --273 ADD R15, R15, R17 //result = result + 4
  when x"00000448" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "100101";  --274 LB, R16, R0,101 //R16 = Mem(101) = 4
  when x"0000044C" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --275 BLT R14, R16, 3
  when x"00000450" => rd <= "000111" & "00000" & "10001" & "00000" & "00001" & "100100";  --276 LB R17, R0, 100 //R17 = Mem(100) = 2 //R17 to hold the amount to be added to result
  when x"00000454" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --277 SUB R14, R14, R16 //a = a - 4
  when x"00000458" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --278 ADD R15, R15, R17 //result = result + 2
  when x"0000045C" => rd <= "000111" & "00000" & "10000" & "00000" & "00001" & "100100";  --279 LB, R16, R0,100 //R16 = Mem(100) = 2
  when x"00000460" => rd <= "001001" & "01110" & "10000" & "00000" & "00000" & "000011";  --280 BLT R14, R16, 3
  when x"00000464" => rd <= "000001" & "00000" & "10001" & "00000" & "00000" & "000001";  --281 ADDI R17, R0, 1 //R17 stores the amount to be added to result
  when x"00000468" => rd <= "000000" & "01110" & "10000" & "01110" & "00000" & "000011";  --282 SUB R14, R14, R16 //a = a - 2
  when x"0000046C" => rd <= "000000" & "01111" & "10001" & "01111" & "00000" & "000001";  --283 ADD R15, R15, R17 //result = result + 1
  when x"00000470" => rd <= "000001" & "01111" & "01110" & "00000" & "00000" & "000000";  --284 ADDI R14, R15, 0 //Store the newly shifted by one value before the next iteration of the loop
  when x"00000474" => rd <= "000001" & "10010" & "10010" & "00000" & "00000" & "000001";  --285 ADDI R18, R18, 1 //R18 increments after each single bit right rotate
  when x"00000478" => rd <= "001010" & "10011" & "10010" & "00000" & "00000" & "000001";  --286 BEQ R18, R19, 1 //If we've shifted right enough times, skip the jump
  when x"0000047C" => rd <= "001100" & "00000" & "00000" & "00000" & "00010" & "000000";  --287 ***CHANGED BY E****JMP 128 //should jump to after the initialization period of the right shift
  when x"00000480" => rd <= "001010" & "00100" & "00000" & "00000" & "00000" & "000101";  --288 BEQ R4, R0, 5
  when x"00000484" => rd <= "001010" & "11011" & "00000" & "00000" & "00000" & "000010";  --289 BEQ R27, R0, 2
  when x"00000488" => rd <= "000010" & "11011" & "11011" & "00000" & "00000" & "000001";  --290 SUBI R27, R27, 1
  when x"0000048C" => rd <= "001100" & "00000" & "00000" & "00000" & "00001" & "110101";  --291 JMP 117
  when x"00000490" => rd <= "000001" & "11011" & "11011" & "00000" & "00000" & "000001";  --292 ADDI R27, R27, 1
  when x"00000494" => rd <= "001100" & "00000" & "00000" & "00000" & "00001" & "100101";  --293 JMP 101
  when x"00000498" => rd <= "001100" & "00000" & "00000" & "00000" & "00000" & "010100";  --294 JMP 20
  when others => rd <= (others => '0');                                                   
end case;                                                                                  
end process;                                                                               
                                                                                           
end rtl;                                                                                                                                                          